class conv_core_output_tr;
    rand int signed out_reg;
endclass
