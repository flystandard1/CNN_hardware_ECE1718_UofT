class dense1_output_tr;
    rand int signed dense_sigmoid[120];
endclass
