class dense2_output_tr;
    rand int dense_sum2[10];
endclass
