class maxpooling_output_tr;
    rand logic signed [15:0] max_layer_out[5][14][14];
endclass
